LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity monitor is
	port
	(

	);
end;

architecture struct of monitor is

begin 

end struct;
