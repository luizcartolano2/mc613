library ieee;
use ieee.std_logic_1164.all;

PACKAGE xbar_v3_package is
	
end xbar_v3_package;
