LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity velha is
	port
	(

	);
end;

architecture struct of velha is

begin 

end struct;
